//////////////////////////////////////////////////////////////////
//  Yusme Pradera ypradera@pdx.edu
//  
// Date: 7/1/2020
//
// testbench for the Behavioral model for a 2^n to n priority encoder.
// 
////////////////////////////////////////////////////////////////
`timescale 1ns/1ps
module designA_netlist_tb();
	// used for # of output bits
  parameter n= 3;
  
     logic [(2**n)-1:0] in;  //2^n bits Input
     logic [n-1:0] out;     //n bits Output 
   
// start stimulus
  initial begin 
    in = 4'b0;
  
    for (int i=0; i < 2**(2**n)-1; i = i+1 ) begin
           #2 in = in + 1'b1;
    end
  end
    
  designA_netlist uut(.in(in),.out(out));
   
  initial begin
    $monitor( "     in=%b :  out=%b    ",in,out);    
   end
  
endmodule
